wire [BW_USERNAME-1:0] username_string = `FORMAT_STRING("None");
wire [BW_GIT_NAME-1:0] home_git_name_string = `FORMAT_STRING("sdk");
wire [BW_GIT_VERSION-1:0] home_git_version_string = `FORMAT_STRING("b43709a");
wire [BW_GIT_VERSION-1:0] devkit_git_version_string = `FORMAT_STRING("cf155e9");
wire [BW_DATE-1:0] design_date_string = `FORMAT_STRING("2026-02-20 18:32");