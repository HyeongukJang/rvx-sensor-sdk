always@(*)
begin : gen_irom_contents
rom_data = 0;
case(rom_index)
0: rom_data = 32'h e1000437;
1: rom_data = 32'h e2011937;
2: rom_data = 32'h 90090913;
3: rom_data = 32'h 00010bb7;
4: rom_data = 32'h 020b8b93;
5: rom_data = 32'h 01740bb3;
6: rom_data = 32'h 000102b7;
7: rom_data = 32'h 00828293;
8: rom_data = 32'h 005402b3;
9: rom_data = 32'h 0002a303;
10: rom_data = 32'h fe030ee3;
11: rom_data = 32'h 000102b7;
12: rom_data = 32'h 005402b3;
13: rom_data = 32'h 0002a303;
14: rom_data = 32'h 00000393;
15: rom_data = 32'h 00730863;
16: rom_data = 32'h 00100393;
17: rom_data = 32'h 02730663;
18: rom_data = 32'h 0240006f;
19: rom_data = 32'h 00200393;
20: rom_data = 32'h 000ba303;
21: rom_data = 32'h fe731ee3;
22: rom_data = 32'h 000102b7;
23: rom_data = 32'h 02828293;
24: rom_data = 32'h 005402b3;
25: rom_data = 32'h 0002a283;
26: rom_data = 32'h 00028067;
27: rom_data = 32'h 0000006f;
28: rom_data = 32'h 000ba303;
29: rom_data = 32'h fc601ce3;
30: rom_data = 32'h 00400393;
31: rom_data = 32'h 00792023;
32: rom_data = 32'h 00300393;
33: rom_data = 32'h 00792223;
34: rom_data = 32'h 000103b7;
35: rom_data = 32'h fff38393;
36: rom_data = 32'h 00792a23;
37: rom_data = 32'h 00200393;
38: rom_data = 32'h 00792c23;
39: rom_data = 32'h 00000393;
40: rom_data = 32'h 00792823;
41: rom_data = 32'h 00100313;
42: rom_data = 32'h 00100393;
43: rom_data = 32'h 007313b3;
44: rom_data = 32'h e2011337;
45: rom_data = 32'h b5030313;
46: rom_data = 32'h 00732023;
47: rom_data = 32'h 000803b7;
48: rom_data = 32'h 04792023;
49: rom_data = 32'h 06092023;
50: rom_data = 32'h 06092223;
51: rom_data = 32'h 06092823;
52: rom_data = 32'h 00100393;
53: rom_data = 32'h 04792823;
54: rom_data = 32'h 04092a23;
55: rom_data = 32'h e10102b7;
56: rom_data = 32'h 08828293;
57: rom_data = 32'h 0002a503;
58: rom_data = 32'h 00350513;
59: rom_data = 32'h 00357293;
60: rom_data = 32'h 40550533;
61: rom_data = 32'h 0d0000ef;
62: rom_data = 32'h 0cc000ef;
63: rom_data = 32'h 0c8000ef;
64: rom_data = 32'h 0c4000ef;
65: rom_data = 32'h 12c000ef;
66: rom_data = 32'h 0a058a63;
67: rom_data = 32'h 00058993;
68: rom_data = 32'h 0b4000ef;
69: rom_data = 32'h 0b0000ef;
70: rom_data = 32'h 0ac000ef;
71: rom_data = 32'h 0a8000ef;
72: rom_data = 32'h 110000ef;
73: rom_data = 32'h 00058a13;
74: rom_data = 32'h 09c000ef;
75: rom_data = 32'h 098000ef;
76: rom_data = 32'h 094000ef;
77: rom_data = 32'h 090000ef;
78: rom_data = 32'h 0f8000ef;
79: rom_data = 32'h 00200313;
80: rom_data = 32'h 02658463;
81: rom_data = 32'h 00400313;
82: rom_data = 32'h 04658463;
83: rom_data = 32'h 00000593;
84: rom_data = 32'h 074000ef;
85: rom_data = 32'h 00ba0023;
86: rom_data = 32'h fff98993;
87: rom_data = 32'h 001a0a13;
88: rom_data = 32'h fe0996e3;
89: rom_data = 32'h f85ff06f;
90: rom_data = 32'h 00000593;
91: rom_data = 32'h 058000ef;
92: rom_data = 32'h 054000ef;
93: rom_data = 32'h 0bc000ef;
94: rom_data = 32'h 0105d593;
95: rom_data = 32'h 00ba1023;
96: rom_data = 32'h ffe98993;
97: rom_data = 32'h 002a0a13;
98: rom_data = 32'h fe0990e3;
99: rom_data = 32'h f5dff06f;
100: rom_data = 32'h 00000593;
101: rom_data = 32'h 030000ef;
102: rom_data = 32'h 02c000ef;
103: rom_data = 32'h 028000ef;
104: rom_data = 32'h 024000ef;
105: rom_data = 32'h 08c000ef;
106: rom_data = 32'h 00ba2023;
107: rom_data = 32'h ffc98993;
108: rom_data = 32'h 004a0a13;
109: rom_data = 32'h fc099ee3;
110: rom_data = 32'h f31ff06f;
111: rom_data = 32'h 000ba023;
112: rom_data = 32'h e8dff06f;
113: rom_data = 32'h 00008b13;
114: rom_data = 32'h 00200393;
115: rom_data = 32'h 00792c23;
116: rom_data = 32'h 000803b7;
117: rom_data = 32'h 00838393;
118: rom_data = 32'h 04792023;
119: rom_data = 32'h 00300613;
120: rom_data = 32'h 088000ef;
121: rom_data = 32'h 01055613;
122: rom_data = 32'h 080000ef;
123: rom_data = 32'h 00855613;
124: rom_data = 32'h 078000ef;
125: rom_data = 32'h 00050613;
126: rom_data = 32'h 070000ef;
127: rom_data = 32'h 000803b7;
128: rom_data = 32'h 04792023;
129: rom_data = 32'h 064000ef;
130: rom_data = 32'h 04c92283;
131: rom_data = 32'h 01f2d313;
132: rom_data = 32'h fe031ce3;
133: rom_data = 32'h 00300393;
134: rom_data = 32'h 00792c23;
135: rom_data = 32'h 00859593;
136: rom_data = 32'h 005585b3;
137: rom_data = 32'h 00150513;
138: rom_data = 32'h 000b0093;
139: rom_data = 32'h 00008067;
140: rom_data = 32'h 0ff00293;
141: rom_data = 32'h 0055f333;
142: rom_data = 32'h 0085d593;
143: rom_data = 32'h 0055f3b3;
144: rom_data = 32'h 0085d593;
145: rom_data = 32'h 0055fe33;
146: rom_data = 32'h 0085d593;
147: rom_data = 32'h 008e1e13;
148: rom_data = 32'h 01c5e5b3;
149: rom_data = 32'h 01039393;
150: rom_data = 32'h 0075e5b3;
151: rom_data = 32'h 01831313;
152: rom_data = 32'h 0065e5b3;
153: rom_data = 32'h 00008067;
154: rom_data = 32'h 04892383;
155: rom_data = 32'h 01f3d393;
156: rom_data = 32'h fe039ce3;
157: rom_data = 32'h 04c92423;
158: rom_data = 32'h 07492383;
159: rom_data = 32'h 0013f393;
160: rom_data = 32'h fe038ce3;
161: rom_data = 32'h 00008067;
endcase
end